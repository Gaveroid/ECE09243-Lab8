module InstMem(addy, inst);

	input [7:0] addy;
	output [31:0] inst;
	
	

endmodule
